`include "q48_0.sv"
`include "q48_1.sv"
`include "q48_tb.sv"
