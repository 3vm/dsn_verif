module tb ;

initial
begin
  $system("grep task *");
end

  logic vikram;
endmodule
