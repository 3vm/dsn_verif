// this is a test module
module mytb; //line comment at end of a line
endmodule
