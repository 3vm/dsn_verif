module tb ;
real p = 0.00513 ;
initial begin
   $display ( "%d" , p ) ;
   $display ( "%f" , p ) ;
   $display ( "%1.2f" , p ) ;
   $display ( "%1.2e" , p ) ;
 end
  logic vikram;
endmodule
