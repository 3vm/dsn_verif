module tb;
  logic p;
  logic q; //wire q;
  
  initial begin
    p = 5;
    //q = 10;
   end
   
   assign q = p;
endmodule