module tb; 
endmodule

/*
Which of these parameter usages is invalid?


Solution
1) port list cannot be modified with generate statement using parameters. 
2) Generate variable names can't be concatenated like in a scripting language like TCL.
3) Generate for loop cannot be inside sensitivity list.
*/