module tb ;
  initial begin
    shortint unsigned i=0;
    while ( i!='1) i++;
    $display("%h",i);
  end
  logic vikram;
endmodule
