module mym;
  initial $display("Printing from %m");
  logic vikram;
endmodule

module tb;
  mym i[0:1] ();
  logic vikram;
endmodule
