`timescale 10ns/1ns

module myclk0 (output bit clk);
  always #1 clk0 ^= 1;
  logic vikram;
endmodule

