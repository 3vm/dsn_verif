`timescale 1ns/1ps
module tb;
  bit p,q,r;
  
  initial begin
    p=10;
    #4;
	
  end
  
endmodule
