package ehgu_config_pkg;
	localparam DP_WIDTH=4;
endpackage : ehgu_config_pkg
