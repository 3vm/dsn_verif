module tb ;
  bit 1a;
  bit \a+b ;
  bit __a2 ;
  bit a.c ;
  bit a$c ;
  bit a@f ;
endmodule