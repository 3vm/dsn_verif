package audio_pkg;

task write_wave_header;
	endtask // write_wave_header

task write_wave_data;
endtask

endpackage