
program tb ;
`include "star.sv"


initial begin
 $display("Song Generated");
 $finish;
end

  logic vikram;
endprogram
