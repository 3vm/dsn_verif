module tb ;
  initial begin
    int k = 2 ** 32 - 1;
    $display ( "%d" , k ) ;
  end
endmodule
