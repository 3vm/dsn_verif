`include "q48_0.sv"
`include "q48_1.sv"
`include "q48_tb.sv"
`include "../thee/thee_clk_freq_meter.sv"
