
module tb ;

timeunit 1ns;
timeprecision 1ps;


initial begin
	$display ( "Hello World" );
end

endmodule
