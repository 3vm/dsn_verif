module tb ;

initial
begin
  $system("grep task *");
end

endmodule
