package chip_config_pkg ;
localparam NUMBUF = 16 ;

localparam NUMREG = 6 ;
localparam BUFEN_ADDR_0 = 0 ;
localparam BUFEN_ADDR_1 = 1 ;
localparam BUFTYPE_ADDR_0 = 2 ;
localparam BUFTYPE_ADDR_1 = 3 ;
localparam ACTDET_ADDR_0 = 4 ;
localparam ACTDET_ADDR_1 = 5 ;
localparam time ACTDET_PERIOD = 100ns ;
endpackage

