
module tb;
byte dmv_customers0;
int dmv_customers1[$];
int dmv_customers2[100];
logic [7:0] dmv_customers3;
  logic vikram;
endmodule