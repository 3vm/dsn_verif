module mym;
  initial $display("Printing from %m");
endmodule

module tb;
  mym i[0:1] ();
endmodule
