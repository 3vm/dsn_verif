continuation of q51
