`timescale 100ps/1ps
