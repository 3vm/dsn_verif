module tb;
  initial begin
    $display("%d",$clog2(3000'd 99999_99999_99999_99999_99999_99999_99999_99999_99999_99999));
    $display("%d",$clog2('d 99999_99999_99999_99999_99999_99999_99999_99999_99999_99999));
  end
endmodule 
