package t ;
endpackage

module tb ;
initial begin
fork
endfork

case ( 0 )
endcase

end

task xyz ;
endtask

  logic vikram;
endmodule
