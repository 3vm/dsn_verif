package thee_mathsci_consts_pkg;
	localparam real const_e=2.71828182846;
	localparam real const_pi=3.14159265359;
//gravitational constant
//mu naught
//epsilon naught

endpackage
