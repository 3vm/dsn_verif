package ehgu_config_pkg;
	localparam DP_WIDTH=16;
endpackage : ehgu_config_pkg
