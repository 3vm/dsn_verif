module mym0
#(parameter N=3)
( input d1, output d2 ,
generate 
  if (N>=3) begin
    input d2, output d3,
  end
endgenerate
 output de
);
endmodule

